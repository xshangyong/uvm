`ifndef GLOBAL_PACKAGE
`define GLOBAL_PACKAGE

package global_package;
	parameter	PACKAGE_DRIVE_NUM = 3;
endpackage

`endif